library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bcd_adder_structural_tb is
-- empty
end bcd_adder_structural_tb;

architecture tb of bcd_adder_structural is
	
begin
end;